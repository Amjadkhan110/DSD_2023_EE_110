module lab4_tb();
 logic [1:0] a1;   
 logic [1:0] b1;
 logic R1;
 logic G1;
 logic B1;
 lab4 UTT(
  .a(a1),
  .b(b1),
  .R(R1),
  .G(G1),
  .B(B1)
);
initial
begin
a1[0]=0;a1[1]=0;b1[0]=0;b1[1]=0;
#10;
a1[0]=0;a1[1]=0;b1[0]=0;b1[1]=1;
#10;
a1[0]=0;a1[1]=0;b1[0]=1;b1[1]=0;
#10;
a1[0]=0;a1[1]=0;b1[0]=1;b1[1]=1;
#10;
a1[0]=0;a1[1]=1;b1[0]=0;b1[1]=0;
#10;
a1[0]=0;a1[1]=1;b1[0]=0;b1[1]=1;
#10;
a1[0]=0;a1[1]=1;b1[0]=1;b1[1]=0;
#10;
a1[0]=0;a1[1]=1;b1[0]=1;b1[1]=1;
#10;
a1[0]=1;a1[1]=0;b1[0]=0;b1[1]=0;
#10;
a1[0]=1;a1[1]=0;b1[0]=0;b1[1]=1;
#10;
a1[0]=1;a1[1]=0;b1[0]=1;b1[1]=0;
#10;
a1[0]=1;a1[1]=0;b1[0]=1;b1[1]=1;
#10;
a1[0]=1;a1[1]=1;b1[0]=0;b1[1]=0;
#10;
a1[0]=1;a1[1]=1;b1[0]=0;b1[1]=1;
#10;
a1[0]=1;a1[1]=1;b1[0]=1;b1[1]=0;
#10;
a1[0]=1;a1[1]=1;b1[0]=1;b1[1]=1;
#10;

$stop;
end
initial
begin
   $monitor("R=%b,G=%b, B_=%b, a[0]=%b,a[1]=%b,b[0]=%b,b[1]=%b", R1,G1,B1,a1[0],a1[1],b1[0],b1[1]);
end
endmodule

